* /home/ameya/esim/eSim-2.0/library/SubcircuitLibrary/swi/swi.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jul 29 12:04:24 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  /d0 /D /gnd /gnd eSim_MOS_N		
M2  /vdd /D /d0 /vdd eSim_MOS_P		
M5  /out /D /vil /vdd eSim_MOS_P		
M3  /out /d0 /vil /gnd eSim_MOS_N		
M6  /vih /D /out /gnd eSim_MOS_N		
M4  /vih /d0 /out /vdd eSim_MOS_P		
U1  /D /vdd /gnd /vil /vih /out PORT		

.end
